module veryl_testcase_Module48;
endmodule

`ifdef __veryl_test_test1__
module test;
   initial begin
       $display("hello");
   end
endmodule

`endif
