module veryl_testcase_Module43;
    StructA          a;
    logic        [10-1:0] b;

    assign b = a.memberA;
endmodule
