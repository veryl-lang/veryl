module veryl_testcase_Module65;
    logic a  ; always_comb a   = 1;
    logic b_n; always_comb b_n = 1;
    logic c  ; always_comb c   = 1;
    logic d  ; always_comb d   = 1;
    logic e  ; always_comb e   = 1;
    logic f  ; always_comb f   = 1;

    logic _x0  ; always_comb _x0   = a;
    logic _x1  ; always_comb _x1   = a;
    logic _x2  ; always_comb _x2   = ~b_n;
    logic _x3  ; always_comb _x3   = b_n;
    logic _x4  ; always_comb _x4   = ~b_n;
    logic _x5  ; always_comb _x5   = b_n;
    logic _x6_n; always_comb _x6_n = ~c;
    logic _x7_n; always_comb _x7_n = d;
    logic _x8_n; always_comb _x8_n = ~e;
    logic _x9_n; always_comb _x9_n = f;
endmodule
//# sourceMappingURL=../map/testcases/sv/65_cast_to_clock_reset.sv.map
