

package veryl_testcase___Package25__1;
    localparam int unsigned C = 1;
    typedef struct packed {
        logic [C-1:0] s;
    } S;
endpackage
//# sourceMappingURL=../map/25_dependency_1.sv.map
