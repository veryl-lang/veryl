module veryl_testcase_Module24;
    (* ram_style="block" *)
    logic _a;
    always_comb _a = 1;
    (* mark_debug="true" *)
    logic _b;
    always_comb _b = 1;
endmodule
