module veryl_testcase_Module62;
    logic clock;
    logic reset;
    logic in   ;
    always_comb in = 0;
    logic out  ;
    always_comb clock = 1;
    always_comb reset = 1;
    always_comb out   = in;
endmodule
//# sourceMappingURL=../map/testcases/sv/62_raw_identifier.sv.map
