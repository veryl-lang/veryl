module veryl_testcase_Module47;
endmodule


module test;
   initial begin
       $display("hello");
   end
endmodule


// comment
