module veryl_testcase_Module24;
    (* ram_style="block" *)
    logic  _a;
    (* mark_debug="true" *)
    logic  _b;
endmodule
