module veryl_testcase_Module22;
    logic     signed [10-1:0] _a;
    always_comb _a = 1;
    tri logic signed [10-1:0] _b;
    assign _b = 1;
    tri logic signed [10-1:0] _c;
    assign _c = 1;
    logic            [10-1:0] _d;
    always_comb _d = 1;
endmodule
//# sourceMappingURL=../map/testcases/sv/22_type_modifier.sv.map
