module veryl_testcase_Module26;
    logic [10-1:0]         _a               ; always_comb _a                = 1;
    logic [10-1:0][10-1:0] _b               ; always_comb _b                = 1;
    logic [10-1:0][10-1:0] _c [0:2-1]       ; always_comb _c = '{1, 1};
    logic [10-1:0][10-1:0] _d [0:2-1][0:2-1]; always_comb _d = '{'{1, 1}, '{1, 1}};
endmodule
//# sourceMappingURL=../map/testcases/sv/26_array.sv.map
