module veryl_testcase_Module34;
    localparam int unsigned a0 = '0;
    localparam int unsigned a1 = '1;
    localparam int unsigned a2 = 'x;
    localparam int unsigned a3 = 'z;
    localparam int unsigned a4 = 10'b0000000000;
    localparam int unsigned a5 = 10'b1111111111;
    localparam int unsigned a6 = 10'bxxxxxxxxxx;
    localparam int unsigned a7 = 10'bzzzzzzzzzz;
endmodule
