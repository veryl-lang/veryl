module Module15 ;
    logic  _a;
    if (1) begin 
    :label
        logic  _a;
    end
    if (1) begin 
    :label1
        logic  _a;
    end
endmodule
