module Module23 #(

    parameter int unsigned ParamA  = 1,
    parameter int unsigned ParamB  = 1,

    parameter int unsigned ParamC  = 1
) (

    input logic  port_a,
    input logic  port_b,

    input logic  port_c
);

    logic [10-1:0] _a;

    logic [10-1:0] _b;logic [10-1:0] _c;

endmodule

module Module23_A;

endmodule

module Module23_B;

endmodulemodule Module23_C;

endmodule
