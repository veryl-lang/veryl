module veryl_testcase_Module33;
    localparam int unsigned a0 = 1'b1;
    localparam int unsigned a1 = 4'b1010;
    localparam int unsigned a2 = 1'o1;
    localparam int unsigned a3 = 10'o1234;
    localparam int unsigned a4 = 1'd1;
    localparam int unsigned a5 = 24'd12345678;
    localparam int unsigned a6 = 1'h1;
    localparam int unsigned a7 = 32'hffffffff;
    localparam int unsigned a8 = 208'hffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff_ffff;
endmodule
//# sourceMappingURL=../map/33_widthless_num.sv.map
