
//# sourceMappingURL=../map/testcases/sv/30_empty.sv.map
