module veryl_testcase_Module57;
    localparam int unsigned     A = veryl_testcase___Package57__1::X;
    localparam longint unsigned B = veryl_testcase___Package57__2::X;
endmodule

package veryl_testcase___Package57__1;
    localparam int unsigned X = 1;
endpackage
package veryl_testcase___Package57__2;
    localparam int unsigned X = 2;
endpackage
