module veryl_testcase_Module22;
    logic     signed [10-1:0] _a;
    tri logic signed [10-1:0] _b;
    tri logic signed [10-1:0] _c;
    logic            [10-1:0] _d;
endmodule
