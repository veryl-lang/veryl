module veryl_testcase_Module26;
    logic [10-1:0]         _a                 ;
    logic [10-1:0][10-1:0] _b                 ;
    logic [10-1:0][10-1:0] _c [0:10-1]        ;
    logic [10-1:0][10-1:0] _d [0:10-1][0:10-1];
endmodule
