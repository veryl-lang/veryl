module veryl_testcase_Module62;
    logic clock;
    logic reset;
    always_comb clock = 1;
    always_comb reset = 1;
endmodule
//# sourceMappingURL=../map/testcases/sv/62_raw_identifier.sv.map
