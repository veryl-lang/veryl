module Module24;
    (* ram_style="block" *)
    logic  _a;
    (* mark_debug="true" *)
    logic  _b;
endmodule
