module veryl_testcase_Module49;
    logic a;

    always_comb begin
        a = $acos();
        a = $acosh();
        a = $asin();
        a = $asinh();
        a = $assertcontrol();
        a = $assertfailoff();
        a = $assertfailon();
        a = $assertkill();
        a = $assertnonvacuouson();
        a = $assertoff();
        a = $asserton();
        a = $assertpassoff();
        a = $assertpasson();
        a = $assertvacuousoff();
        a = $async$and$array();
        a = $async$and$plane();
        a = $async$nand$array();
        a = $async$nand$plane();
        a = $async$nor$array();
        a = $async$nor$plane();
        a = $async$or$array();
        a = $async$or$plane();
        a = $atan();
        a = $atan2();
        a = $atanh();
        a = $bits(logic);
        a = $bitstoreal();
        a = $bitstoshortreal();
        a = $cast();
        a = $ceil();
        a = $changed();
        a = $changed_gclk();
        a = $changing_gclk();
        a = $clog2(1);
        a = $cos();
        a = $cosh();
        a = $countbits();
        a = $countones();
        a = $coverage_control();
        a = $coverage_get();
        a = $coverage_get_max();
        a = $coverage_merge();
        a = $coverage_save();
        a = $dimensions();
        a = $display();
        a = $displayb();
        a = $displayh();
        a = $displayo();
        a = $dist_chi_square();
        a = $dist_erlang();
        a = $dist_exponential();
        a = $dist_normal();
        a = $dist_poisson();
        a = $dist_t();
        a = $dist_uniform();
        a = $dumpall();
        a = $dumpfile();
        a = $dumpflush();
        a = $dumplimit();
        a = $dumpoff();
        a = $dumpon();
        a = $dumpports();
        a = $dumpportsall();
        a = $dumpportsflush();
        a = $dumpportslimit();
        a = $dumpportsoff();
        a = $dumpportson();
        a = $dumpvars();
        a = $error();
        a = $exit();
        a = $exp();
        a = $falling_gclk();
        a = $fatal();
        a = $fclose();
        a = $fdisplay();
        a = $fdisplayb();
        a = $fdisplayh();
        a = $fdisplayo();
        a = $fell();
        a = $fell_gclk();
        a = $feof();
        a = $ferror();
        a = $fflush();
        a = $fgetc();
        a = $fgets();
        a = $finish();
        a = $floor();
        a = $fmonitor();
        a = $fmonitorb();
        a = $fmonitorh();
        a = $fmonitoro();
        a = $fopen();
        a = $fread();
        a = $fscanf();
        a = $fseek();
        a = $fstrobe();
        a = $fstrobeb();
        a = $fstrobeh();
        a = $fstrobeo();
        a = $ftell();
        a = $future_gclk();
        a = $fwrite();
        a = $fwriteb();
        a = $fwriteh();
        a = $fwriteo();
        a = $get_coverage();
        a = $high();
        a = $hypot();
        a = $increment();
        a = $info();
        a = $isunbounded();
        a = $isunknown();
        a = $itor();
        a = $left();
        a = $ln();
        a = $load_coverage_db();
        a = $log10();
        a = $low();
        a = $monitor();
        a = $monitorb();
        a = $monitorh();
        a = $monitoro();
        a = $monitoroff();
        a = $monitoron();
        a = $onehot();
        a = $onehot0();
        a = $past();
        a = $past_gclk();
        a = $pow();
        a = $printtimescale();
        a = $q_add();
        a = $q_exam();
        a = $q_full();
        a = $q_initialize();
        a = $q_remove();
        a = $random();
        a = $readmemb();
        a = $readmemh();
        a = $realtime();
        a = $realtobits();
        a = $rewind();
        a = $right();
        a = $rising_gclk();
        a = $rose();
        a = $rose_gclk();
        a = $rtoi();
        a = $sampled();
        a = $set_coverage_db_name();
        a = $sformat();
        a = $sformatf();
        a = $shortrealtobits();
        a = $signed();
        a = $sin();
        a = $sinh();
        a = $size();
        a = $sqrt();
        a = $sscanf();
        a = $stable();
        a = $stable_gclk();
        a = $steady_gclk();
        a = $stime();
        a = $stop();
        a = $strobe();
        a = $strobeb();
        a = $strobeh();
        a = $strobeo();
        a = $swrite();
        a = $swriteb();
        a = $swriteh();
        a = $swriteo();
        a = $sync$and$array();
        a = $sync$and$plane();
        a = $sync$nand$array();
        a = $sync$nand$plane();
        a = $sync$nor$array();
        a = $sync$nor$plane();
        a = $sync$or$array();
        a = $sync$or$plane();
        a = $system();
        a = $tan();
        a = $tanh();
        a = $test$plusargs();
        a = $time();
        a = $timeformat();
        a = $typename();
        a = $ungetc();
        a = $unpacked_dimensions();
        a = $unsigned();
        a = $value$plusargs();
        a = $warning();
        a = $write();
        a = $writeb();
        a = $writeh();
        a = $writememb();
        a = $writememh();
        a = $writeo();
    end
endmodule

package veryl_testcase_Package49;
    localparam int unsigned a = 1;
    localparam int unsigned b = $clog2(a);
endpackage
//# sourceMappingURL=../map/49_system_function.sv.map
