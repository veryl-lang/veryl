module veryl_testcase_Module52;
endmodule
module test;
   initial begin
       $display("hello");
   end
endmodule

