module veryl_testcase_Module27;
    localparam string a = "aaa";

    string _b;
    always_comb _b = "bbb";
endmodule
