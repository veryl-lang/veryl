


module veryl_testcase_Module69A #(
    parameter int unsigned A = 1,
    parameter int unsigned B = 1,
    parameter int unsigned C = 1
) (
    input  var logic a,
    input  var logic b,
    output var logic c
);
    always_comb c = a;
endmodule
//# sourceMappingURL=../map/69_proto.sv.map
