module veryl_testcase_Module34;
    logic [32-1:0] _a0; always_comb _a0 = '0;
    logic [32-1:0] _a1; always_comb _a1 = '1;
    logic [32-1:0] _a2; always_comb _a2 = 'x;
    logic [32-1:0] _a3; always_comb _a3 = 'z;
    logic [32-1:0] _a4; always_comb _a4 = 10'b0000000000;
    logic [32-1:0] _a5; always_comb _a5 = 10'b1111111111;
    logic [32-1:0] _a6; always_comb _a6 = 10'bxxxxxxxxxx;
    logic [32-1:0] _a7; always_comb _a7 = 10'bzzzzzzzzzz;
endmodule
//# sourceMappingURL=../map/testcases/sv/34_width_all_set.sv.map
