
//# sourceMappingURL=../map/30_empty.sv.map
