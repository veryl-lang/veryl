package veryl_testcase_Package59A;
    localparam int unsigned XLEN = 32;
endpackage

package veryl_testcase_Package59B;
    localparam int unsigned XLEN = veryl_testcase_Package59A::XLEN;
endpackage
