module veryl_testcase_Module68;
    std_fifo u (
        .i_clk         (),
        .i_rst         (),
        .i_clear       (),
        .o_empty       (),
        .o_almost_full (),
        .o_full        (),
        .o_word_count  (),
        .i_push        (),
        .i_data        (),
        .i_pop         (),
        .o_data        ()
    );
endmodule
//# sourceMappingURL=../map/testcases/sv/68_std.sv.map
