module veryl_testcase_Module27;
    localparam string a = "aaa";

    string _b;
    assign _b = "bbb";
endmodule
