module Module15 ;
    logic  a;
    if (1) begin :label
        logic  a;
    end
    if (1) begin :label1
        logic  a;
    end
endmodule
