module veryl_testcase_Module31;
    initial begin
        $display("initial");
    end

    final begin
        $display("final");
    end
endmodule
