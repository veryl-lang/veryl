


module veryl_testcase_Module19
    import PackageA::A;
    import PackageA::*;
;
    import PackageA::A;
    import PackageA::*;
endmodule

interface veryl_testcase_Interface19
    import PackageA::A;
    import PackageA::*;
;
    import PackageA::A;
    import PackageA::*;
endinterface

package veryl_testcase_Package19;
    import PackageA::A;
    import PackageA::*;
    import PackageA::A;
    import PackageA::*;
    export PackageA::A;
    export *::*;
endpackage
