module veryl_testcase_Module37;
    int unsigned _a;
    assign _a = veryl_testcase_Package37::A;
endmodule
package veryl_testcase_Package37;
    localparam int unsigned A = 1;
endpackage
