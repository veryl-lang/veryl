



module veryl_testcase_Module25A
    import veryl_sample4___bar_pkg__32::*;
    import veryl_sample4___baz_pkg__veryl_testcase___Package25__1_C::*;
(
    input var logic                    i_clk  ,
    input var logic                    i_rst_n,
    veryl_sample3_data_if.mp_in  in_if  ,
    veryl_sample3_data_if.mp_out out_if 
);



    veryl_sample3_data_if data_if ();

    veryl_sample_delay u0 (
        .i_clk     (i_clk       ),
        .i_rst_n_n (i_rst_n     ),
        .i_d       (in_if.data  ),
        .o_d       (data_if.data)
    );

    veryl_sample2_delay u1 (
        .i_clk     (i_clk       ),
        .i_rst_n_n (i_rst_n     ),
        .i_d       (data_if.data),
        .o_d       (out_if.data )
    );

    veryl_sample4___bar_module__veryl_sample4___foo_pkg__veryl_sample4___bar_pkg__32_BAR__veryl_sample4___bar_pkg__32 u2 ();
endmodule

module veryl_testcase___Module25B____Package25__1;
    import veryl_testcase___Package25__1::*;


    veryl_sample4___qux_if__veryl_testcase___Package25__1_S u3       ();
    veryl_sample4___qux_if__veryl_testcase___Package25__1_S u4       ();
    always_comb u3.qux.s = '0;
    always_comb u4.qux.s = '0;
endmodule

module veryl_testcase_Module25C;
    veryl_testcase___Module25B____Package25__1 u5 ();
endmodule
//# sourceMappingURL=../map/25_dependency_2.sv.map
