module veryl_testcase_Module43;
    StructA          a;
    logic   [10-1:0] b;

    always_comb b = a.memberA;
endmodule
//# sourceMappingURL=../map/testcases/sv/43_sv_member.sv.map
