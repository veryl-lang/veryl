


module veryl_testcase_Module69A #(
    parameter int unsigned A = 1,
    parameter int unsigned B = 1,
    parameter int unsigned C = 1
) (
    input  logic a,
    input  logic b,
    output logic c
);
    always_comb c = a;
endmodule
//# sourceMappingURL=../map/testcases/sv/69_proto.sv.map
