module veryl_testcase_Module22;
    logic     signed [10-1:0] _a;
    always_comb _a = 1;
    tri logic signed [10-1:0] _b;
    always_comb _b = 1;
    tri logic signed [10-1:0] _c;
    always_comb _c = 1;
    logic            [10-1:0] _d;
    always_comb _d = 1;
endmodule
