module veryl_testcase_Module31;
    initial begin
        $display("initial");
    end

    final begin
        $display("final");
    end
endmodule
//# sourceMappingURL=../map/testcases/sv/31_initial_final.sv.map
